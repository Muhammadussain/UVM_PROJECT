///////////////////////////////////////////////////////////////////////////////
// File:        cfs_apb_types.sv
// Author:      Cristian Florin Slav
// Date:        2023-07-05
// Description: Types used by the APB agent
///////////////////////////////////////////////////////////////////////////////
`ifndef CFS_APB_TYPES_SV
  `define CFS_APB_TYPES_SV

    //Virtual interface type
    typedef virtual cfs_apb_if cfs_apb_vif;

`endif